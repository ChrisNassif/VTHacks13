
module bridge (
	clk_clk,
	memory_mem_a,
	memory_mem_ba,
	memory_mem_ck,
	memory_mem_ck_n,
	memory_mem_cke,
	memory_mem_cs_n,
	memory_mem_ras_n,
	memory_mem_cas_n,
	memory_mem_we_n,
	memory_mem_reset_n,
	memory_mem_dq,
	memory_mem_dqs,
	memory_mem_dqs_n,
	memory_mem_odt,
	memory_mem_dm,
	memory_oct_rzqin,
	hps_io_hps_io_usb0_inst_D0,
	hps_io_hps_io_usb0_inst_D1,
	hps_io_hps_io_usb0_inst_D2,
	hps_io_hps_io_usb0_inst_D3,
	hps_io_hps_io_usb0_inst_D4,
	hps_io_hps_io_usb0_inst_D5,
	hps_io_hps_io_usb0_inst_D6,
	hps_io_hps_io_usb0_inst_D7,
	hps_io_hps_io_usb0_inst_CLK,
	hps_io_hps_io_usb0_inst_STP,
	hps_io_hps_io_usb0_inst_DIR,
	hps_io_hps_io_usb0_inst_NXT,
	button_external_export);	

	input		clk_clk;
	output	[12:0]	memory_mem_a;
	output	[2:0]	memory_mem_ba;
	output		memory_mem_ck;
	output		memory_mem_ck_n;
	output		memory_mem_cke;
	output		memory_mem_cs_n;
	output		memory_mem_ras_n;
	output		memory_mem_cas_n;
	output		memory_mem_we_n;
	output		memory_mem_reset_n;
	inout	[7:0]	memory_mem_dq;
	inout		memory_mem_dqs;
	inout		memory_mem_dqs_n;
	output		memory_mem_odt;
	output		memory_mem_dm;
	input		memory_oct_rzqin;
	inout		hps_io_hps_io_usb0_inst_D0;
	inout		hps_io_hps_io_usb0_inst_D1;
	inout		hps_io_hps_io_usb0_inst_D2;
	inout		hps_io_hps_io_usb0_inst_D3;
	inout		hps_io_hps_io_usb0_inst_D4;
	inout		hps_io_hps_io_usb0_inst_D5;
	inout		hps_io_hps_io_usb0_inst_D6;
	inout		hps_io_hps_io_usb0_inst_D7;
	input		hps_io_hps_io_usb0_inst_CLK;
	output		hps_io_hps_io_usb0_inst_STP;
	input		hps_io_hps_io_usb0_inst_DIR;
	input		hps_io_hps_io_usb0_inst_NXT;
	input		button_external_export;
endmodule
