// (C) 2001-2024 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files from any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel FPGA IP License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
// agreement for further details.


module uart_small_hps_0_hps_io_border(
// memory
  output wire [13 - 1 : 0 ] mem_a
 ,output wire [3 - 1 : 0 ] mem_ba
 ,output wire [1 - 1 : 0 ] mem_ck
 ,output wire [1 - 1 : 0 ] mem_ck_n
 ,output wire [1 - 1 : 0 ] mem_cke
 ,output wire [1 - 1 : 0 ] mem_cs_n
 ,output wire [1 - 1 : 0 ] mem_ras_n
 ,output wire [1 - 1 : 0 ] mem_cas_n
 ,output wire [1 - 1 : 0 ] mem_we_n
 ,output wire [1 - 1 : 0 ] mem_reset_n
 ,inout wire [8 - 1 : 0 ] mem_dq
 ,inout wire [1 - 1 : 0 ] mem_dqs
 ,inout wire [1 - 1 : 0 ] mem_dqs_n
 ,output wire [1 - 1 : 0 ] mem_odt
 ,output wire [1 - 1 : 0 ] mem_dm
 ,input wire [1 - 1 : 0 ] oct_rzqin
// hps_io
 ,inout wire [1 - 1 : 0 ] hps_io_usb0_inst_D0
 ,inout wire [1 - 1 : 0 ] hps_io_usb0_inst_D1
 ,inout wire [1 - 1 : 0 ] hps_io_usb0_inst_D2
 ,inout wire [1 - 1 : 0 ] hps_io_usb0_inst_D3
 ,inout wire [1 - 1 : 0 ] hps_io_usb0_inst_D4
 ,inout wire [1 - 1 : 0 ] hps_io_usb0_inst_D5
 ,inout wire [1 - 1 : 0 ] hps_io_usb0_inst_D6
 ,inout wire [1 - 1 : 0 ] hps_io_usb0_inst_D7
 ,input wire [1 - 1 : 0 ] hps_io_usb0_inst_CLK
 ,output wire [1 - 1 : 0 ] hps_io_usb0_inst_STP
 ,input wire [1 - 1 : 0 ] hps_io_usb0_inst_DIR
 ,input wire [1 - 1 : 0 ] hps_io_usb0_inst_NXT
);

assign hps_io_usb0_inst_D0 = intermediate[1] ? intermediate[0] : 'z;
assign hps_io_usb0_inst_D1 = intermediate[3] ? intermediate[2] : 'z;
assign hps_io_usb0_inst_D2 = intermediate[5] ? intermediate[4] : 'z;
assign hps_io_usb0_inst_D3 = intermediate[7] ? intermediate[6] : 'z;
assign hps_io_usb0_inst_D4 = intermediate[9] ? intermediate[8] : 'z;
assign hps_io_usb0_inst_D5 = intermediate[11] ? intermediate[10] : 'z;
assign hps_io_usb0_inst_D6 = intermediate[13] ? intermediate[12] : 'z;
assign hps_io_usb0_inst_D7 = intermediate[15] ? intermediate[14] : 'z;

wire [16 - 1 : 0] intermediate;

cyclonev_hps_peripheral_usb usb0_inst(
 .USB_ULPI_STP({
    hps_io_usb0_inst_STP[0:0] // 0:0
  })
,.USB_ULPI_DATA_I({
    hps_io_usb0_inst_D7[0:0] // 7:7
   ,hps_io_usb0_inst_D6[0:0] // 6:6
   ,hps_io_usb0_inst_D5[0:0] // 5:5
   ,hps_io_usb0_inst_D4[0:0] // 4:4
   ,hps_io_usb0_inst_D3[0:0] // 3:3
   ,hps_io_usb0_inst_D2[0:0] // 2:2
   ,hps_io_usb0_inst_D1[0:0] // 1:1
   ,hps_io_usb0_inst_D0[0:0] // 0:0
  })
,.USB_ULPI_NXT({
    hps_io_usb0_inst_NXT[0:0] // 0:0
  })
,.USB_ULPI_DIR({
    hps_io_usb0_inst_DIR[0:0] // 0:0
  })
,.USB_ULPI_DATA_O({
    intermediate[14:14] // 7:7
   ,intermediate[12:12] // 6:6
   ,intermediate[10:10] // 5:5
   ,intermediate[8:8] // 4:4
   ,intermediate[6:6] // 3:3
   ,intermediate[4:4] // 2:2
   ,intermediate[2:2] // 1:1
   ,intermediate[0:0] // 0:0
  })
,.USB_ULPI_CLK({
    hps_io_usb0_inst_CLK[0:0] // 0:0
  })
,.USB_ULPI_DATA_OE({
    intermediate[15:15] // 7:7
   ,intermediate[13:13] // 6:6
   ,intermediate[11:11] // 5:5
   ,intermediate[9:9] // 4:4
   ,intermediate[7:7] // 3:3
   ,intermediate[5:5] // 2:2
   ,intermediate[3:3] // 1:1
   ,intermediate[1:1] // 0:0
  })
);


hps_sdram hps_sdram_inst(
 .mem_dq({
    mem_dq[7:0] // 7:0
  })
,.mem_odt({
    mem_odt[0:0] // 0:0
  })
,.mem_ras_n({
    mem_ras_n[0:0] // 0:0
  })
,.mem_dqs_n({
    mem_dqs_n[0:0] // 0:0
  })
,.mem_dqs({
    mem_dqs[0:0] // 0:0
  })
,.mem_dm({
    mem_dm[0:0] // 0:0
  })
,.mem_we_n({
    mem_we_n[0:0] // 0:0
  })
,.mem_cas_n({
    mem_cas_n[0:0] // 0:0
  })
,.mem_ba({
    mem_ba[2:0] // 2:0
  })
,.mem_a({
    mem_a[12:0] // 12:0
  })
,.mem_cs_n({
    mem_cs_n[0:0] // 0:0
  })
,.mem_ck({
    mem_ck[0:0] // 0:0
  })
,.mem_cke({
    mem_cke[0:0] // 0:0
  })
,.oct_rzqin({
    oct_rzqin[0:0] // 0:0
  })
,.mem_reset_n({
    mem_reset_n[0:0] // 0:0
  })
,.mem_ck_n({
    mem_ck_n[0:0] // 0:0
  })
);

endmodule

