module array_uart_transmitter #(
    parameter CLOCK_FREQ = 50_000_000,
    parameter BAUD_RATE = 115200
)(
    input wire clk,
    input wire rst_n,
    input wire [31:0] data_array,
    input wire send_trigger,        // Pulse to start transmission
    output wire uart_tx,
    output wire busy
);

    // UART transmitter signals
    wire [7:0] tx_data;
    wire tx_valid;
    wire tx_ready;
    
    // State machine for array transmission
    typedef enum logic [2:0] {
        IDLE,
        TRANSMIT_HEADER,
        TRANSMIT_DATA,
        TRANSMIT_FOOTER
    } state_t;
    
    state_t state;
    reg [3:0] array_index;
    reg [1:0] byte_index;
    reg [31:0] current_word;
    
    // UART transmitter instance
    uart_tx #(
        .CLOCK_FREQ(CLOCK_FREQ),
        .BAUD_RATE(BAUD_RATE)
    ) uart_transmitter (
        .clk(clk),
        .rst_n(rst_n),
        .data(tx_data),
        .valid(tx_valid),
        .ready(tx_ready),
        .tx(uart_tx)
    );
    
    // Control logic
    reg send_trigger_prev;
    wire send_edge;
    
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            send_trigger_prev <= 1'b0;
        end else begin
            send_trigger_prev <= send_trigger;
        end
    end
    
    assign send_edge = send_trigger && !send_trigger_prev;
    assign busy = (state != IDLE);
    
    // Transmission state machine
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state <= IDLE;
            array_index <= 0;
            byte_index <= 0;
            current_word <= 32'h00000000;
        end else begin
            case (state)
                IDLE: begin
                    if (send_edge) begin
                        state <= TRANSMIT_HEADER;
                        array_index <= 0;
                        byte_index <= 0;
                    end
                end
                
                TRANSMIT_HEADER: begin
                    if (tx_valid && tx_ready) begin
                        state <= TRANSMIT_DATA;
                        current_word <= data_array[0];
                        array_index <= 0;
                        byte_index <= 0;
                    end
                end
                
                TRANSMIT_DATA: begin
                    if (tx_valid && tx_ready) begin
                        if (byte_index == 3) begin
                            // Finished current word
                            if (array_index == 0) begin
                                // Finished all words
                                state <= TRANSMIT_FOOTER;
                            end else begin
                                // Move to next word
                                array_index <= array_index + 1;
                                current_word <= data_array[array_index + 1];
                                byte_index <= 0;
                            end
                        end else begin
                            // Move to next byte
                            byte_index <= byte_index + 1;
                        end
                    end
                end
                
                TRANSMIT_FOOTER: begin
                    if (tx_valid && tx_ready) begin
                        state <= IDLE;
                    end
                end
            endcase
        end
    end
    
    // Data multiplexer
    reg [7:0] tx_data_reg;
    reg tx_valid_reg;
    
    always_comb begin
        case (state)
            TRANSMIT_HEADER: begin
                tx_data_reg = 8'hAA;  // Header byte
                tx_valid_reg = 1'b1;
            end
            
            TRANSMIT_DATA: begin
                case (byte_index)
                    2'b00: tx_data_reg = current_word[7:0];
                    2'b01: tx_data_reg = current_word[15:8];
                    2'b10: tx_data_reg = current_word[23:16];
                    2'b11: tx_data_reg = current_word[31:24];
                endcase
                tx_valid_reg = 1'b1;
            end
            
            TRANSMIT_FOOTER: begin
                tx_data_reg = 8'h55;  // Footer byte
                tx_valid_reg = 1'b1;
            end
            
            default: begin
                tx_data_reg = 8'h00;
                tx_valid_reg = 1'b0;
            end
        endcase
    end
    
    assign tx_data = tx_data_reg;
    assign tx_valid = tx_valid_reg;

endmodule